library verilog;
use verilog.vl_types.all;
entity test_bench3 is
    generic(
        n               : integer := 2
    );
end test_bench3;
