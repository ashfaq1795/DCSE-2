library verilog;
use verilog.vl_types.all;
entity test_bench4 is
end test_bench4;
