library verilog;
use verilog.vl_types.all;
entity tb_buffer is
end tb_buffer;
