library verilog;
use verilog.vl_types.all;
entity stim_mux8x1 is
end stim_mux8x1;
