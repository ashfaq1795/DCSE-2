library verilog;
use verilog.vl_types.all;
entity stim_mux2x1 is
end stim_mux2x1;
