library verilog;
use verilog.vl_types.all;
entity stimdec3x8 is
end stimdec3x8;
