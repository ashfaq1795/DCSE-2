library verilog;
use verilog.vl_types.all;
entity stimmux2x1 is
end stimmux2x1;
