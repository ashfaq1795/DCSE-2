module carry(c,A,B);
input A,B;
output c;
assign c=A&B;
endmodule
