library verilog;
use verilog.vl_types.all;
entity stimmux4x1 is
end stimmux4x1;
