library verilog;
use verilog.vl_types.all;
entity stim_mux4x1 is
end stim_mux4x1;
