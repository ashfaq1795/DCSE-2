library verilog;
use verilog.vl_types.all;
entity stim_half_sub is
end stim_half_sub;
