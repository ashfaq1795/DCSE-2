library verilog;
use verilog.vl_types.all;
entity stim_adder is
end stim_adder;
