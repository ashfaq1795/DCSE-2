library verilog;
use verilog.vl_types.all;
entity test_bench2 is
    generic(
        n               : integer := 2
    );
end test_bench2;
