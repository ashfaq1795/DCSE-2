library verilog;
use verilog.vl_types.all;
entity test_bench3 is
end test_bench3;
