library verilog;
use verilog.vl_types.all;
entity stimdecode is
end stimdecode;
