library verilog;
use verilog.vl_types.all;
entity test_4_bits_adder is
end test_4_bits_adder;
