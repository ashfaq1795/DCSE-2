library verilog;
use verilog.vl_types.all;
entity stim_d is
end stim_d;
