module CARRY (C, A, B);
 
	output C;
	input A, B;
	
	and a1 (C, A, B);
	
endmodule