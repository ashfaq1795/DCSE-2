library verilog;
use verilog.vl_types.all;
entity test_bench4 is
    generic(
        n               : integer := 7
    );
end test_bench4;
