library verilog;
use verilog.vl_types.all;
entity stimg1 is
end stimg1;
