library verilog;
use verilog.vl_types.all;
entity stimdec2x4 is
end stimdec2x4;
