library verilog;
use verilog.vl_types.all;
entity test_bench2 is
end test_bench2;
