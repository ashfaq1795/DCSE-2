library verilog;
use verilog.vl_types.all;
entity test_bench1 is
end test_bench1;
