library verilog;
use verilog.vl_types.all;
entity equation is
    port(
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        x4              : in     vl_logic;
        x5              : in     vl_logic;
        z               : out    vl_logic
    );
end equation;
